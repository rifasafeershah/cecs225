// Code your design here
module adder4bit(
  input [3:0] A,B,
  output [3:0] SUM
);
  assign SUM = A + B;
endmodule
